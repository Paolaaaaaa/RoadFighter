///*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module SC_STATEMACHINE #(parameter MUX41_SELECTWIDTH=32)(
	//////////// OUTPUTS //////////
	
	SC_STATEMACHINE_SIGNAL_OUT,
	
	SC_STATEMACHINE_SIGNAL_OUT_1,
	SC_STATEMACHINE_SIGNAL_OUT_2,
	SC_STATEMACHINE_SIGNAL_OUT_3,
	SC_STATEMACHINE_SIGNAL_OUT_4,
	SC_STATEMACHINE_SIGNAL_OUT_5,
	SC_STATEMACHINE_SIGNAL_OUT_6,
	SC_STATEMACHINE_SIGNAL_OUT_7,
	//////////// INPUTS //////////
	SC_STATEMACHINE_CONTADOR_T,
	SC_STATEMACHINE_RESET_INHigh,
	SC_STATEMACHINE_START_INLow,
	SC_STATEMACHONE_CLOCK_50,
	SC_STATEMACHINE_COMPARATOR,
	SC_STATEMACHINE_CONTADOR_LV
);	
//=======================================================
//  PARAMETER declarations
//=========
//=============================================

output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_Timer;

output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_1_Timer_cte;
output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_2_Load;
output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_3_MUX_SEL_1;
output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_4_MUX_SEL_2;
output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_5_MUX_SEL_3;
//output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_6;
//output	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_7;


input  	SC_STATEMACHINE_CONTADOR_T;
input 	SC_STATEMACHINE_RESET_INHigh;
input 	SC_STATEMACHINE_START_INLow;
input		SC_STATEMACHINE_CLOCK_50;
input		SC_STATEMACHINE_COMPARATOR;
input 	SC_STATEMACHINE_CONTADOR_LV;

reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_reg;

reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_1_reg;
reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_2_reg;
reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_3_reg;
reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_4_reg;
reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_5_reg;
//reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_6_reg;
//reg	[MUX41_SELECTWIDTH-1:0]  SC_STATEMACHINE_SIGNAL_OUT_7_reg;

reg	[MUX41_SELECTWIDTH-1:0] SC_TATEMACHINE_CTE_reg_1;
reg	[MUX41_SELECTWIDTH-1:0] SC_STATEMACHINE_CTE_reg_2;

reg	[MUX41_SELECTWIDTH-1:0] SC_STATEMACHINE_CTE_reg_3;
reg	[MUX41_SELECTWIDTH-1:0] SC_STATEMACHINE_CTE_reg_4;

reg	[MUX41_SELECTWIDTH-1:0] SC_STATEMACHINE_CTE_reg_5;
reg	[MUX41_SELECTWIDTH-1:0] SC_STATEMACHINE_CTE_reg_6;


always @(*)
begin
   if(SC_STATEMACHINE_CONTADOR_LV <=8'b000001010)// LV hasta 10, cada 0.35s genera un load
		SC_STATEMACHINE_SIGNAL_OUT_reg = SC_STATEMACHINE_CLOCK_50_reg;
		SC_STATEMACHINE_SIGNAL_OUT_1_reg = 32'b00000001000010110000011101100000*SC_STATEMACHINE_CTE_reg_1;
		
	else if(SC_STATEMACHINE_CONTADOR_LV >=8'b000001010 && SC_STATEMACHINE_CONTADOR_LV<=8'b00010001)
		SC_STATEMACHINE_SIGNAL_OUT_3_reg = 1b'1;
	
	else if (SC_STATEMACHINE_CONTADOR_LV >=8'b00010001 && SC_STATEMACHINE_CONTADOR_LV<=8'b000100000)//LV 11 hasta 32, cada 0.3s genera un load
		SC_STATEMACHINE_SIGNAL_OUT_reg = SC_STATEMACHINE_CLOCK_50;
		SC_STATEMACHINE_SIGNAL_OUT_1_reg = 32'b00000000111001001110000111000000*SC_STATEMACHINE_CTE_reg_3;
		
	else if(SC_STATEMACHINE_CONTADOR_LV >=8'b000100000 && SC_STATEMACHINE_CONTADOR_LV<=8'b00100111)
		SC_STATEMACHINE_SIGNAL_OUT_4_reg = 1b'1;
		
	else if (SC_STATEMACHINE_CONTADOR_LV >=8'b00100111 && SC_STATEMACHINE_CONTADOR_LV<=8'b00111011)//LV 11 hasta 32, cada 0.3s genera un load
		SC_STATEMACHINE_SIGNAL_OUT_reg = SC_STATEMACHINE_CLOCK_50;
		SC_STATEMACHINE_SIGNAL_OUT_1_reg = 32'b00000000101111101011110000100000*SC_STATEMACHINE_CTE_reg_5;
		
	else
		SC_STATEMACHINE_SIGNAL_OUT_reg = 32'b00000000000000000000000000000000;
		
//   else if( SC_STATEMACHINE_RESET_INHigh == 1 && SC_STATEMACHINE_CONTADOR  == 1)/// cuando reset == 1 pantalla en 0 unos
//   begin   	
//	  SC_STATEMACHINE_SIGNAL_OUT_1_reg= 0;
//
//	  SC_STATEMACHINE_SIGNAL_OUT_2_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_3_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_4_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_5_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_6_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_7_reg= 0;
//	  SC_STATEMACHINE_SIGNAL_OUT_reg= 0;
//	end	
//   else // está en 2 saca el random
//	begin	
//	  SC_STATEMACHINE_SIGNAL_OUT_1_reg= 2;
//
//	  SC_STATEMACHINE_SIGNAL_OUT_2_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_3_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_4_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_5_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_6_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_7_reg= 2;
//	  SC_STATEMACHINE_SIGNAL_OUT_reg= 2;
//		
//	end

end

begin
	if (SC_STATEMACHINE_CONTADOR_T == 1'b1)
		SC_STATEMACHINE_SIGNAL_OUT_2_reg = 1b'1
		SC_STATEMACHINE_SIGNAL_OUT_5_reg = 1b'1
	else 
		SC_STATEMACHINE_SIGNAL_OUT_2_Load = 1b'0
		SC_STATEMACHINE_SIGNAL_OUT_5_reg = 1b'0
		
end


assign SC_STATEMACHINE_SIGNAL_OUT_Timer = SC_STATEMACHINE_SIGNAL_OUT_reg;

assign SC_STATEMACHINE_SIGNAL_OUT_1_Timer_cte = SC_STATEMACHINE_SIGNAL_OUT_1_reg;
assign SC_STATEMACHINE_SIGNAL_OUT_2_Load = SC_STATEMACHINE_SIGNAL_OUT_2_reg;
assign SC_STATEMACHINE_SIGNAL_OUT_3_MUX_SEL_1 = SC_STATEMACHINE_SIGNAL_OUT_3_reg;
assign SC_STATEMACHINE_SIGNAL_OUT_4_MUX_SEL_2 = SC_STATEMACHINE_SIGNAL_OUT_4_reg;
assign SC_STATEMACHINE_SIGNAL_OUT_5_MUX_SEL_3 = SC_STATEMACHINE_SIGNAL_OUT_5_reg;

assign SC_TATEMACHINE_CTE_reg_1 = SC_STATEMACHINE_CTE_reg_2+25'b0000000000000000000000001;
assign SC_STATEMACHINE_CTE_reg_2 = SC_TATEMACHINE_CTE_reg_1;

assign SC_TATEMACHINE_CTE_reg_3 = SC_STATEMACHINE_CTE_reg_4+25'b0000000000000000000000001;
assign SC_STATEMACHINE_CTE_reg_4 = SC_TATEMACHINE_CTE_reg_3;

assign SC_TATEMACHINE_CTE_reg_5 = SC_STATEMACHINE_CTE_reg_6+25'b0000000000000000000000001;
assign SC_STATEMACHINE_CTE_reg_6 = SC_TATEMACHINE_CTE_reg_5;


//assign SC_STATEMACHINE_SIGNAL_OUT_1 = SC_STATEMACHINE_SIGNAL_OUT_1_reg;
//
//assign  SC_STATEMACHINE_SIGNAL_OUT_2 = SC_STATEMACHINE_SIGNAL_OUT_2_reg;
//assign  SC_STATEMACHINE_SIGNAL_OUT_3 = SC_STATEMACHINE_SIGNAL_OUT_3_reg;
//assign SC_STATEMACHINE_SIGNAL_OUT_4 = SC_STATEMACHINE_SIGNAL_OUT_4_reg;
//assign SC_STATEMACHINE_SIGNAL_OUT_5 = SC_STATEMACHINE_SIGNAL_OUT_5_reg;
//assign SC_STATEMACHINE_SIGNAL_OUT_6 = SC_STATEMACHINE_SIGNAL_OUT_6_reg;
//assign SC_STATEMACHINE_SIGNAL_OUT_7 =SC_STATEMACHINE_SIGNAL_OUT_7_reg;
//assign SC_STATEMACHINE_SIGNAL_OUT = SC_STATEMACHINE_SIGNAL_OUT_reg;

 
 endmodule
